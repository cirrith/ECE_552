/********************************************************************************************************
/		MODULE: Fetch
/		PURPOSE: First pipeline section of processor, get instruction from instruction memory
/
/		INPUTS: clk -
				rst_n - 
				
/				
/		OUTPUTS: 
********************************************************************************************************/
module Fetch();

Instruction memory

endmodule