/****************************
purpose: Given a 16 bit input perform the given opcode by 8 when sh is high
****************************/

module shift8 (in, op, sh, out);
input [15:0] in;
input sh;
input [1:0] op;

output out;






endmodule 
