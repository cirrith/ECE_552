moudle ALU_tb.sv