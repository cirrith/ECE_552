module ShRL(In, Amt, Out);

// Declare inputs and outputs
input [3:0] Amt;
input [15:0] In;
output [15:0] Out;

// Declare wires



////////////////////////////////////////////////////////////////////////////////
////////////////////		 	Do the thing!				////////////////////
////////////////////////////////////////////////////////////////////////////////




endmodule