module PC_inc(Curr_PC, Inc_PC);

	input [15:0] Curr_PC;

	output [15:0] Inc_PC;

	assign Inc_PC = ;

endmodule