/****************************
purpose: Given a 16 bit input perform the given opcode by 2 when sh is high
****************************/

module shift2 (in, op, sh, out);
input [15:0] in;
input sh;
input [1:0] op;

output out;






endmodule 
