/********************************************************************************************************
/		MODULE: Execute
/		PURPOSE: Given all the possible inputs to the alu and the corresponding control signals perform
/				the command.
/
/		INPUTS: 
/
/		OUTPUTS: 
********************************************************************************************************/
module Execute();

ALU

endmodule