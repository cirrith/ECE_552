module mux4x4_1(A, B, C, D, Sel, Out);

// Declare inputs and outputs
input [15:0] A, B, C, D;
input [1:0] Sel;
output [15:0] Out;


////////////////////////////////////////////////////////////////////////////////
////////////////////		 	Do the thing!				////////////////////
////////////////////////////////////////////////////////////////////////////////


mux4_1 multi_mux[15:0](.A(A), .B(B), .C(C), .D(D), .Sel(Sel), .Out(Out));


endmodule