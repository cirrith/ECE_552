/********************************************************************************************************
/		MODULE: Decode
/		PURPOSE: Contain the control and register_file 
/
/		INPUTS: 
/
/		OUTPUTS: 
********************************************************************************************************/
module Decode();

Register File
Register File Input
Extender
Control

endmodule