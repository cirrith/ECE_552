library verilog;
use verilog.vl_types.all;
entity proc_hier_pbench is
end proc_hier_pbench;
